module smcauth(clk, rst, g_input, e_input, o);
  input clk;
  input [255:0] e_input;
  input [255:0] g_input;
  output o;
  input rst;
  wire W1;
  wire W2;
  wire W3;
  wire W4;
  wire W5;
  wire W6;
  wire W7;
  wire W8;
  wire W9;
  wire W10;
  wire W11;
  wire W12;
  wire W13;
  wire W14;
  wire W15;
  wire W16;
  wire W17;
  wire W18;
  wire W19;
  wire W20;
  wire W21;
  wire W22;
  wire W23;
  wire W24;
  wire W25;
  wire W26;
  wire W27;
  wire W28;
  wire W29;
  wire W30;
  wire W31;
  wire W32;
  wire W33;
  wire W34;
  wire W35;
  wire W36;
  wire W37;
  wire W38;
  wire W39;
  wire W40;
  wire W41;
  wire W42;
  wire W43;
  wire W44;
  wire W45;
  wire W46;
  wire W47;
  wire W48;
  wire W49;
  wire W50;
  wire W51;
  wire W52;
  wire W53;
  wire W54;
  wire W55;
  wire W56;
  wire W57;
  wire W58;
  wire W59;
  wire W60;
  wire W61;
  wire W62;
  wire W63;
  wire W64;
  wire W65;
  wire W66;
  wire W67;
  wire W68;
  wire W69;
  wire W70;
  wire W71;
  wire W72;
  wire W73;
  wire W74;
  wire W75;
  wire W76;
  wire W77;
  wire W78;
  wire W79;
  wire W80;
  wire W81;
  wire W82;
  wire W83;
  wire W84;
  wire W85;
  wire W86;
  wire W87;
  wire W88;
  wire W89;
  wire W90;
  wire W91;
  wire W92;
  wire W93;
  wire W94;
  wire W95;
  wire W96;
  wire W97;
  wire W98;
  wire W99;
  wire W100;
  wire W101;
  wire W102;
  wire W103;
  wire W104;
  wire W105;
  wire W106;
  wire W107;
  wire W108;
  wire W109;
  wire W110;
  wire W111;
  wire W112;
  wire W113;
  wire W114;
  wire W115;
  wire W116;
  wire W117;
  wire W118;
  wire W119;
  wire W120;
  wire W121;
  wire W122;
  wire W123;
  wire W124;
  wire W125;
  wire W126;
  wire W127;
  wire W128;
  wire W129;
  wire W130;
  wire W131;
  wire W132;
  wire W133;
  wire W134;
  wire W135;
  wire W136;
  wire W137;
  wire W138;
  wire W139;
  wire W140;
  wire W141;
  wire W142;
  wire W143;
  wire W144;
  wire W145;
  wire W146;
  wire W147;
  wire W148;
  wire W149;
  wire W150;
  wire W151;
  wire W152;
  wire W153;
  wire W154;
  wire W155;
  wire W156;
  wire W157;
  wire W158;
  wire W159;
  wire W160;
  wire W161;
  wire W162;
  wire W163;
  wire W164;
  wire W165;
  wire W166;
  wire W167;
  wire W168;
  wire W169;
  wire W170;
  wire W171;
  wire W172;
  wire W173;
  wire W174;
  wire W175;
  wire W176;
  wire W177;
  wire W178;
  wire W179;
  wire W180;
  wire W181;
  wire W182;
  wire W183;
  wire W184;
  wire W185;
  wire W186;
  wire W187;
  wire W188;
  wire W189;
  wire W190;
  wire W191;
  wire W192;
  wire W193;
  wire W194;
  wire W195;
  wire W196;
  wire W197;
  wire W198;
  wire W199;
  wire W200;
  wire W201;
  wire W202;
  wire W203;
  wire W204;
  wire W205;
  wire W206;
  wire W207;
  wire W208;
  wire W209;
  wire W210;
  wire W211;
  wire W212;
  wire W213;
  wire W214;
  wire W215;
  wire W216;
  wire W217;
  wire W218;
  wire W219;
  wire W220;
  wire W221;
  wire W222;
  wire W223;
  wire W224;
  wire W225;
  wire W226;
  wire W227;
  wire W228;
  wire W229;
  wire W230;
  wire W231;
  wire W232;
  wire W233;
  wire W234;
  wire W235;
  wire W236;
  wire W237;
  wire W238;
  wire W239;
  wire W240;
  wire W241;
  wire W242;
  wire W243;
  wire W244;
  wire W245;
  wire W246;
  wire W247;
  wire W248;
  wire W249;
  wire W250;
  wire W251;
  wire W252;
  wire W253;
  wire W254;
  wire W255;
  wire W256;
  wire W257;
  wire W258;
  wire W259;
  wire W260;
  wire W261;
  wire W262;
  wire W263;
  wire W264;
  wire W265;
  wire W266;
  wire W267;
  wire W268;
  wire W269;
  wire W270;
  wire W271;
  wire W272;
  wire W273;
  wire W274;
  wire W275;
  wire W276;
  wire W277;
  wire W278;
  wire W279;
  wire W280;
  wire W281;
  wire W282;
  wire W283;
  wire W284;
  wire W285;
  wire W286;
  wire W287;
  wire W288;
  wire W289;
  wire W290;
  wire W291;
  wire W292;
  wire W293;
  wire W294;
  wire W295;
  wire W296;
  wire W297;
  wire W298;
  wire W299;
  wire W300;
  wire W301;
  wire W302;
  wire W303;
  wire W304;
  wire W305;
  wire W306;
  wire W307;
  wire W308;
  wire W309;
  wire W310;
  wire W311;
  wire W312;
  wire W313;
  wire W314;
  wire W315;
  wire W316;
  wire W317;
  wire W318;
  wire W319;
  wire W320;
  wire W321;
  wire W322;
  wire W323;
  wire W324;
  wire W325;
  wire W326;
  wire W327;
  wire W328;
  wire W329;
  wire W330;
  wire W331;
  wire W332;
  wire W333;
  wire W334;
  wire W335;
  wire W336;
  wire W337;
  wire W338;
  wire W339;
  wire W340;
  wire W341;
  wire W342;
  wire W343;
  wire W344;
  wire W345;
  wire W346;
  wire W347;
  wire W348;
  wire W349;
  wire W350;
  wire W351;
  wire W352;
  wire W353;
  wire W354;
  wire W355;
  wire W356;
  wire W357;
  wire W358;
  wire W359;
  wire W360;
  wire W361;
  wire W362;
  wire W363;
  wire W364;
  wire W365;
  wire W366;
  wire W367;
  wire W368;
  wire W369;
  wire W370;
  wire W371;
  wire W372;
  wire W373;
  wire W374;
  wire W375;
  wire W376;
  wire W377;
  wire W378;
  wire W379;
  wire W380;
  wire W381;
  wire W382;
  wire W383;
  wire W384;
  wire W385;
  wire W386;
  wire W387;
  wire W388;
  wire W389;
  wire W390;
  wire W391;
  wire W392;
  wire W393;
  wire W394;
  wire W395;
  wire W396;
  wire W397;
  wire W398;
  wire W399;
  wire W400;
  wire W401;
  wire W402;
  wire W403;
  wire W404;
  wire W405;
  wire W406;
  wire W407;
  wire W408;
  wire W409;
  wire W410;
  wire W411;
  wire W412;
  wire W413;
  wire W414;
  wire W415;
  wire W416;
  wire W417;
  wire W418;
  wire W419;
  wire W420;
  wire W421;
  wire W422;
  wire W423;
  wire W424;
  wire W425;
  wire W426;
  wire W427;
  wire W428;
  wire W429;
  wire W430;
  wire W431;
  wire W432;
  wire W433;
  wire W434;
  wire W435;
  wire W436;
  wire W437;
  wire W438;
  wire W439;
  wire W440;
  wire W441;
  wire W442;
  wire W443;
  wire W444;
  wire W445;
  wire W446;
  wire W447;
  wire W448;
  wire W449;
  wire W450;
  wire W451;
  wire W452;
  wire W453;
  wire W454;
  wire W455;
  wire W456;
  wire W457;
  wire W458;
  wire W459;
  wire W460;
  wire W461;
  wire W462;
  wire W463;
  wire W464;
  wire W465;
  wire W466;
  wire W467;
  wire W468;
  wire W469;
  wire W470;
  wire W471;
  wire W472;
  wire W473;
  wire W474;
  wire W475;
  wire W476;
  wire W477;
  wire W478;
  wire W479;
  wire W480;
  wire W481;
  wire W482;
  wire W483;
  wire W484;
  wire W485;
  wire W486;
  wire W487;
  wire W488;
  wire W489;
  wire W490;
  wire W491;
  wire W492;
  wire W493;
  wire W494;
  wire W495;
  wire W496;
  wire W497;
  wire W498;
  wire W499;
  wire W500;
  wire W501;
  wire W502;
  wire W503;
  wire W504;
  wire W505;
  wire W506;
  wire W507;
  wire W508;
  wire W509;
  wire W510;

  OR C1 (
    .A(g_input[0]),
    .B(e_input[0]),
    .Z(W1)
  );

  OR C2 (
    .A(g_input[1]),
    .B(W1),
    .Z(W2)
  );

  OR C3 (
    .A(e_input[1]),
    .B(W2),
    .Z(W3)
  );

  OR C4 (
    .A(g_input[2]),
    .B(W3),
    .Z(W4)
  );

  OR C5 (
    .A(e_input[2]),
    .B(W4),
    .Z(W5)
  );

  OR C6 (
    .A(g_input[3]),
    .B(W5),
    .Z(W6)
  );

  OR C7 (
    .A(e_input[3]),
    .B(W6),
    .Z(W7)
  );

  OR C8 (
    .A(g_input[4]),
    .B(W7),
    .Z(W8)
  );

  OR C9 (
    .A(e_input[4]),
    .B(W8),
    .Z(W9)
  );

  OR C10 (
    .A(g_input[5]),
    .B(W9),
    .Z(W10)
  );

  OR C11 (
    .A(e_input[5]),
    .B(W10),
    .Z(W11)
  );

  OR C12 (
    .A(g_input[6]),
    .B(W11),
    .Z(W12)
  );

  OR C13 (
    .A(e_input[6]),
    .B(W12),
    .Z(W13)
  );

  OR C14 (
    .A(g_input[7]),
    .B(W13),
    .Z(W14)
  );

  OR C15 (
    .A(e_input[7]),
    .B(W14),
    .Z(W15)
  );

  OR C16 (
    .A(g_input[8]),
    .B(W15),
    .Z(W16)
  );

  OR C17 (
    .A(e_input[8]),
    .B(W16),
    .Z(W17)
  );

  OR C18 (
    .A(g_input[9]),
    .B(W17),
    .Z(W18)
  );

  OR C19 (
    .A(e_input[9]),
    .B(W18),
    .Z(W19)
  );

  OR C20 (
    .A(g_input[10]),
    .B(W19),
    .Z(W20)
  );

  OR C21 (
    .A(e_input[10]),
    .B(W20),
    .Z(W21)
  );

  OR C22 (
    .A(g_input[11]),
    .B(W21),
    .Z(W22)
  );

  OR C23 (
    .A(e_input[11]),
    .B(W22),
    .Z(W23)
  );

  OR C24 (
    .A(g_input[12]),
    .B(W23),
    .Z(W24)
  );

  OR C25 (
    .A(e_input[12]),
    .B(W24),
    .Z(W25)
  );

  OR C26 (
    .A(g_input[13]),
    .B(W25),
    .Z(W26)
  );

  OR C27 (
    .A(e_input[13]),
    .B(W26),
    .Z(W27)
  );

  OR C28 (
    .A(g_input[14]),
    .B(W27),
    .Z(W28)
  );

  OR C29 (
    .A(e_input[14]),
    .B(W28),
    .Z(W29)
  );

  OR C30 (
    .A(g_input[15]),
    .B(W29),
    .Z(W30)
  );

  OR C31 (
    .A(e_input[15]),
    .B(W30),
    .Z(W31)
  );

  OR C32 (
    .A(g_input[16]),
    .B(W31),
    .Z(W32)
  );

  OR C33 (
    .A(e_input[16]),
    .B(W32),
    .Z(W33)
  );

  OR C34 (
    .A(g_input[17]),
    .B(W33),
    .Z(W34)
  );

  OR C35 (
    .A(e_input[17]),
    .B(W34),
    .Z(W35)
  );

  OR C36 (
    .A(g_input[18]),
    .B(W35),
    .Z(W36)
  );

  OR C37 (
    .A(e_input[18]),
    .B(W36),
    .Z(W37)
  );

  OR C38 (
    .A(g_input[19]),
    .B(W37),
    .Z(W38)
  );

  OR C39 (
    .A(e_input[19]),
    .B(W38),
    .Z(W39)
  );

  OR C40 (
    .A(g_input[20]),
    .B(W39),
    .Z(W40)
  );

  OR C41 (
    .A(e_input[20]),
    .B(W40),
    .Z(W41)
  );

  OR C42 (
    .A(g_input[21]),
    .B(W41),
    .Z(W42)
  );

  OR C43 (
    .A(e_input[21]),
    .B(W42),
    .Z(W43)
  );

  OR C44 (
    .A(g_input[22]),
    .B(W43),
    .Z(W44)
  );

  OR C45 (
    .A(e_input[22]),
    .B(W44),
    .Z(W45)
  );

  OR C46 (
    .A(g_input[23]),
    .B(W45),
    .Z(W46)
  );

  OR C47 (
    .A(e_input[23]),
    .B(W46),
    .Z(W47)
  );

  OR C48 (
    .A(g_input[24]),
    .B(W47),
    .Z(W48)
  );

  OR C49 (
    .A(e_input[24]),
    .B(W48),
    .Z(W49)
  );

  OR C50 (
    .A(g_input[25]),
    .B(W49),
    .Z(W50)
  );

  OR C51 (
    .A(e_input[25]),
    .B(W50),
    .Z(W51)
  );

  OR C52 (
    .A(g_input[26]),
    .B(W51),
    .Z(W52)
  );

  OR C53 (
    .A(e_input[26]),
    .B(W52),
    .Z(W53)
  );

  OR C54 (
    .A(g_input[27]),
    .B(W53),
    .Z(W54)
  );

  OR C55 (
    .A(e_input[27]),
    .B(W54),
    .Z(W55)
  );

  OR C56 (
    .A(g_input[28]),
    .B(W55),
    .Z(W56)
  );

  OR C57 (
    .A(e_input[28]),
    .B(W56),
    .Z(W57)
  );

  OR C58 (
    .A(g_input[29]),
    .B(W57),
    .Z(W58)
  );

  OR C59 (
    .A(e_input[29]),
    .B(W58),
    .Z(W59)
  );

  OR C60 (
    .A(g_input[30]),
    .B(W59),
    .Z(W60)
  );

  OR C61 (
    .A(e_input[30]),
    .B(W60),
    .Z(W61)
  );

  OR C62 (
    .A(g_input[31]),
    .B(W61),
    .Z(W62)
  );

  OR C63 (
    .A(e_input[31]),
    .B(W62),
    .Z(W63)
  );

  OR C64 (
    .A(g_input[32]),
    .B(W63),
    .Z(W64)
  );

  OR C65 (
    .A(e_input[32]),
    .B(W64),
    .Z(W65)
  );

  OR C66 (
    .A(g_input[33]),
    .B(W65),
    .Z(W66)
  );

  OR C67 (
    .A(e_input[33]),
    .B(W66),
    .Z(W67)
  );

  OR C68 (
    .A(g_input[34]),
    .B(W67),
    .Z(W68)
  );

  OR C69 (
    .A(e_input[34]),
    .B(W68),
    .Z(W69)
  );

  OR C70 (
    .A(g_input[35]),
    .B(W69),
    .Z(W70)
  );

  OR C71 (
    .A(e_input[35]),
    .B(W70),
    .Z(W71)
  );

  OR C72 (
    .A(g_input[36]),
    .B(W71),
    .Z(W72)
  );

  OR C73 (
    .A(e_input[36]),
    .B(W72),
    .Z(W73)
  );

  OR C74 (
    .A(g_input[37]),
    .B(W73),
    .Z(W74)
  );

  OR C75 (
    .A(e_input[37]),
    .B(W74),
    .Z(W75)
  );

  OR C76 (
    .A(g_input[38]),
    .B(W75),
    .Z(W76)
  );

  OR C77 (
    .A(e_input[38]),
    .B(W76),
    .Z(W77)
  );

  OR C78 (
    .A(g_input[39]),
    .B(W77),
    .Z(W78)
  );

  OR C79 (
    .A(e_input[39]),
    .B(W78),
    .Z(W79)
  );

  OR C80 (
    .A(g_input[40]),
    .B(W79),
    .Z(W80)
  );

  OR C81 (
    .A(e_input[40]),
    .B(W80),
    .Z(W81)
  );

  OR C82 (
    .A(g_input[41]),
    .B(W81),
    .Z(W82)
  );

  OR C83 (
    .A(e_input[41]),
    .B(W82),
    .Z(W83)
  );

  OR C84 (
    .A(g_input[42]),
    .B(W83),
    .Z(W84)
  );

  OR C85 (
    .A(e_input[42]),
    .B(W84),
    .Z(W85)
  );

  OR C86 (
    .A(g_input[43]),
    .B(W85),
    .Z(W86)
  );

  OR C87 (
    .A(e_input[43]),
    .B(W86),
    .Z(W87)
  );

  OR C88 (
    .A(g_input[44]),
    .B(W87),
    .Z(W88)
  );

  OR C89 (
    .A(e_input[44]),
    .B(W88),
    .Z(W89)
  );

  OR C90 (
    .A(g_input[45]),
    .B(W89),
    .Z(W90)
  );

  OR C91 (
    .A(e_input[45]),
    .B(W90),
    .Z(W91)
  );

  OR C92 (
    .A(g_input[46]),
    .B(W91),
    .Z(W92)
  );

  OR C93 (
    .A(e_input[46]),
    .B(W92),
    .Z(W93)
  );

  OR C94 (
    .A(g_input[47]),
    .B(W93),
    .Z(W94)
  );

  OR C95 (
    .A(e_input[47]),
    .B(W94),
    .Z(W95)
  );

  OR C96 (
    .A(g_input[48]),
    .B(W95),
    .Z(W96)
  );

  OR C97 (
    .A(e_input[48]),
    .B(W96),
    .Z(W97)
  );

  OR C98 (
    .A(g_input[49]),
    .B(W97),
    .Z(W98)
  );

  OR C99 (
    .A(e_input[49]),
    .B(W98),
    .Z(W99)
  );

  OR C100 (
    .A(g_input[50]),
    .B(W99),
    .Z(W100)
  );

  OR C101 (
    .A(e_input[50]),
    .B(W100),
    .Z(W101)
  );

  OR C102 (
    .A(g_input[51]),
    .B(W101),
    .Z(W102)
  );

  OR C103 (
    .A(e_input[51]),
    .B(W102),
    .Z(W103)
  );

  OR C104 (
    .A(g_input[52]),
    .B(W103),
    .Z(W104)
  );

  OR C105 (
    .A(e_input[52]),
    .B(W104),
    .Z(W105)
  );

  OR C106 (
    .A(g_input[53]),
    .B(W105),
    .Z(W106)
  );

  OR C107 (
    .A(e_input[53]),
    .B(W106),
    .Z(W107)
  );

  OR C108 (
    .A(g_input[54]),
    .B(W107),
    .Z(W108)
  );

  OR C109 (
    .A(e_input[54]),
    .B(W108),
    .Z(W109)
  );

  OR C110 (
    .A(g_input[55]),
    .B(W109),
    .Z(W110)
  );

  OR C111 (
    .A(e_input[55]),
    .B(W110),
    .Z(W111)
  );

  OR C112 (
    .A(g_input[56]),
    .B(W111),
    .Z(W112)
  );

  OR C113 (
    .A(e_input[56]),
    .B(W112),
    .Z(W113)
  );

  OR C114 (
    .A(g_input[57]),
    .B(W113),
    .Z(W114)
  );

  OR C115 (
    .A(e_input[57]),
    .B(W114),
    .Z(W115)
  );

  OR C116 (
    .A(g_input[58]),
    .B(W115),
    .Z(W116)
  );

  OR C117 (
    .A(e_input[58]),
    .B(W116),
    .Z(W117)
  );

  OR C118 (
    .A(g_input[59]),
    .B(W117),
    .Z(W118)
  );

  OR C119 (
    .A(e_input[59]),
    .B(W118),
    .Z(W119)
  );

  OR C120 (
    .A(g_input[60]),
    .B(W119),
    .Z(W120)
  );

  OR C121 (
    .A(e_input[60]),
    .B(W120),
    .Z(W121)
  );

  OR C122 (
    .A(g_input[61]),
    .B(W121),
    .Z(W122)
  );

  OR C123 (
    .A(e_input[61]),
    .B(W122),
    .Z(W123)
  );

  OR C124 (
    .A(g_input[62]),
    .B(W123),
    .Z(W124)
  );

  OR C125 (
    .A(e_input[62]),
    .B(W124),
    .Z(W125)
  );

  OR C126 (
    .A(g_input[63]),
    .B(W125),
    .Z(W126)
  );

  OR C127 (
    .A(e_input[63]),
    .B(W126),
    .Z(W127)
  );

  OR C128 (
    .A(g_input[64]),
    .B(W127),
    .Z(W128)
  );

  OR C129 (
    .A(e_input[64]),
    .B(W128),
    .Z(W129)
  );

  OR C130 (
    .A(g_input[65]),
    .B(W129),
    .Z(W130)
  );

  OR C131 (
    .A(e_input[65]),
    .B(W130),
    .Z(W131)
  );

  OR C132 (
    .A(g_input[66]),
    .B(W131),
    .Z(W132)
  );

  OR C133 (
    .A(e_input[66]),
    .B(W132),
    .Z(W133)
  );

  OR C134 (
    .A(g_input[67]),
    .B(W133),
    .Z(W134)
  );

  OR C135 (
    .A(e_input[67]),
    .B(W134),
    .Z(W135)
  );

  OR C136 (
    .A(g_input[68]),
    .B(W135),
    .Z(W136)
  );

  OR C137 (
    .A(e_input[68]),
    .B(W136),
    .Z(W137)
  );

  OR C138 (
    .A(g_input[69]),
    .B(W137),
    .Z(W138)
  );

  OR C139 (
    .A(e_input[69]),
    .B(W138),
    .Z(W139)
  );

  OR C140 (
    .A(g_input[70]),
    .B(W139),
    .Z(W140)
  );

  OR C141 (
    .A(e_input[70]),
    .B(W140),
    .Z(W141)
  );

  OR C142 (
    .A(g_input[71]),
    .B(W141),
    .Z(W142)
  );

  OR C143 (
    .A(e_input[71]),
    .B(W142),
    .Z(W143)
  );

  OR C144 (
    .A(g_input[72]),
    .B(W143),
    .Z(W144)
  );

  OR C145 (
    .A(e_input[72]),
    .B(W144),
    .Z(W145)
  );

  OR C146 (
    .A(g_input[73]),
    .B(W145),
    .Z(W146)
  );

  OR C147 (
    .A(e_input[73]),
    .B(W146),
    .Z(W147)
  );

  OR C148 (
    .A(g_input[74]),
    .B(W147),
    .Z(W148)
  );

  OR C149 (
    .A(e_input[74]),
    .B(W148),
    .Z(W149)
  );

  OR C150 (
    .A(g_input[75]),
    .B(W149),
    .Z(W150)
  );

  OR C151 (
    .A(e_input[75]),
    .B(W150),
    .Z(W151)
  );

  OR C152 (
    .A(g_input[76]),
    .B(W151),
    .Z(W152)
  );

  OR C153 (
    .A(e_input[76]),
    .B(W152),
    .Z(W153)
  );

  OR C154 (
    .A(g_input[77]),
    .B(W153),
    .Z(W154)
  );

  OR C155 (
    .A(e_input[77]),
    .B(W154),
    .Z(W155)
  );

  OR C156 (
    .A(g_input[78]),
    .B(W155),
    .Z(W156)
  );

  OR C157 (
    .A(e_input[78]),
    .B(W156),
    .Z(W157)
  );

  OR C158 (
    .A(g_input[79]),
    .B(W157),
    .Z(W158)
  );

  OR C159 (
    .A(e_input[79]),
    .B(W158),
    .Z(W159)
  );

  OR C160 (
    .A(g_input[80]),
    .B(W159),
    .Z(W160)
  );

  OR C161 (
    .A(e_input[80]),
    .B(W160),
    .Z(W161)
  );

  OR C162 (
    .A(g_input[81]),
    .B(W161),
    .Z(W162)
  );

  OR C163 (
    .A(e_input[81]),
    .B(W162),
    .Z(W163)
  );

  OR C164 (
    .A(g_input[82]),
    .B(W163),
    .Z(W164)
  );

  OR C165 (
    .A(e_input[82]),
    .B(W164),
    .Z(W165)
  );

  OR C166 (
    .A(g_input[83]),
    .B(W165),
    .Z(W166)
  );

  OR C167 (
    .A(e_input[83]),
    .B(W166),
    .Z(W167)
  );

  OR C168 (
    .A(g_input[84]),
    .B(W167),
    .Z(W168)
  );

  OR C169 (
    .A(e_input[84]),
    .B(W168),
    .Z(W169)
  );

  OR C170 (
    .A(g_input[85]),
    .B(W169),
    .Z(W170)
  );

  OR C171 (
    .A(e_input[85]),
    .B(W170),
    .Z(W171)
  );

  OR C172 (
    .A(g_input[86]),
    .B(W171),
    .Z(W172)
  );

  OR C173 (
    .A(e_input[86]),
    .B(W172),
    .Z(W173)
  );

  OR C174 (
    .A(g_input[87]),
    .B(W173),
    .Z(W174)
  );

  OR C175 (
    .A(e_input[87]),
    .B(W174),
    .Z(W175)
  );

  OR C176 (
    .A(g_input[88]),
    .B(W175),
    .Z(W176)
  );

  OR C177 (
    .A(e_input[88]),
    .B(W176),
    .Z(W177)
  );

  OR C178 (
    .A(g_input[89]),
    .B(W177),
    .Z(W178)
  );

  OR C179 (
    .A(e_input[89]),
    .B(W178),
    .Z(W179)
  );

  OR C180 (
    .A(g_input[90]),
    .B(W179),
    .Z(W180)
  );

  OR C181 (
    .A(e_input[90]),
    .B(W180),
    .Z(W181)
  );

  OR C182 (
    .A(g_input[91]),
    .B(W181),
    .Z(W182)
  );

  OR C183 (
    .A(e_input[91]),
    .B(W182),
    .Z(W183)
  );

  OR C184 (
    .A(g_input[92]),
    .B(W183),
    .Z(W184)
  );

  OR C185 (
    .A(e_input[92]),
    .B(W184),
    .Z(W185)
  );

  OR C186 (
    .A(g_input[93]),
    .B(W185),
    .Z(W186)
  );

  OR C187 (
    .A(e_input[93]),
    .B(W186),
    .Z(W187)
  );

  OR C188 (
    .A(g_input[94]),
    .B(W187),
    .Z(W188)
  );

  OR C189 (
    .A(e_input[94]),
    .B(W188),
    .Z(W189)
  );

  OR C190 (
    .A(g_input[95]),
    .B(W189),
    .Z(W190)
  );

  OR C191 (
    .A(e_input[95]),
    .B(W190),
    .Z(W191)
  );

  OR C192 (
    .A(g_input[96]),
    .B(W191),
    .Z(W192)
  );

  OR C193 (
    .A(e_input[96]),
    .B(W192),
    .Z(W193)
  );

  OR C194 (
    .A(g_input[97]),
    .B(W193),
    .Z(W194)
  );

  OR C195 (
    .A(e_input[97]),
    .B(W194),
    .Z(W195)
  );

  OR C196 (
    .A(g_input[98]),
    .B(W195),
    .Z(W196)
  );

  OR C197 (
    .A(e_input[98]),
    .B(W196),
    .Z(W197)
  );

  OR C198 (
    .A(g_input[99]),
    .B(W197),
    .Z(W198)
  );

  OR C199 (
    .A(e_input[99]),
    .B(W198),
    .Z(W199)
  );

  OR C200 (
    .A(g_input[100]),
    .B(W199),
    .Z(W200)
  );

  OR C201 (
    .A(e_input[100]),
    .B(W200),
    .Z(W201)
  );

  OR C202 (
    .A(g_input[101]),
    .B(W201),
    .Z(W202)
  );

  OR C203 (
    .A(e_input[101]),
    .B(W202),
    .Z(W203)
  );

  OR C204 (
    .A(g_input[102]),
    .B(W203),
    .Z(W204)
  );

  OR C205 (
    .A(e_input[102]),
    .B(W204),
    .Z(W205)
  );

  OR C206 (
    .A(g_input[103]),
    .B(W205),
    .Z(W206)
  );

  OR C207 (
    .A(e_input[103]),
    .B(W206),
    .Z(W207)
  );

  OR C208 (
    .A(g_input[104]),
    .B(W207),
    .Z(W208)
  );

  OR C209 (
    .A(e_input[104]),
    .B(W208),
    .Z(W209)
  );

  OR C210 (
    .A(g_input[105]),
    .B(W209),
    .Z(W210)
  );

  OR C211 (
    .A(e_input[105]),
    .B(W210),
    .Z(W211)
  );

  OR C212 (
    .A(g_input[106]),
    .B(W211),
    .Z(W212)
  );

  OR C213 (
    .A(e_input[106]),
    .B(W212),
    .Z(W213)
  );

  OR C214 (
    .A(g_input[107]),
    .B(W213),
    .Z(W214)
  );

  OR C215 (
    .A(e_input[107]),
    .B(W214),
    .Z(W215)
  );

  OR C216 (
    .A(g_input[108]),
    .B(W215),
    .Z(W216)
  );

  OR C217 (
    .A(e_input[108]),
    .B(W216),
    .Z(W217)
  );

  OR C218 (
    .A(g_input[109]),
    .B(W217),
    .Z(W218)
  );

  OR C219 (
    .A(e_input[109]),
    .B(W218),
    .Z(W219)
  );

  OR C220 (
    .A(g_input[110]),
    .B(W219),
    .Z(W220)
  );

  OR C221 (
    .A(e_input[110]),
    .B(W220),
    .Z(W221)
  );

  OR C222 (
    .A(g_input[111]),
    .B(W221),
    .Z(W222)
  );

  OR C223 (
    .A(e_input[111]),
    .B(W222),
    .Z(W223)
  );

  OR C224 (
    .A(g_input[112]),
    .B(W223),
    .Z(W224)
  );

  OR C225 (
    .A(e_input[112]),
    .B(W224),
    .Z(W225)
  );

  OR C226 (
    .A(g_input[113]),
    .B(W225),
    .Z(W226)
  );

  OR C227 (
    .A(e_input[113]),
    .B(W226),
    .Z(W227)
  );

  OR C228 (
    .A(g_input[114]),
    .B(W227),
    .Z(W228)
  );

  OR C229 (
    .A(e_input[114]),
    .B(W228),
    .Z(W229)
  );

  OR C230 (
    .A(g_input[115]),
    .B(W229),
    .Z(W230)
  );

  OR C231 (
    .A(e_input[115]),
    .B(W230),
    .Z(W231)
  );

  OR C232 (
    .A(g_input[116]),
    .B(W231),
    .Z(W232)
  );

  OR C233 (
    .A(e_input[116]),
    .B(W232),
    .Z(W233)
  );

  OR C234 (
    .A(g_input[117]),
    .B(W233),
    .Z(W234)
  );

  OR C235 (
    .A(e_input[117]),
    .B(W234),
    .Z(W235)
  );

  OR C236 (
    .A(g_input[118]),
    .B(W235),
    .Z(W236)
  );

  OR C237 (
    .A(e_input[118]),
    .B(W236),
    .Z(W237)
  );

  OR C238 (
    .A(g_input[119]),
    .B(W237),
    .Z(W238)
  );

  OR C239 (
    .A(e_input[119]),
    .B(W238),
    .Z(W239)
  );

  OR C240 (
    .A(g_input[120]),
    .B(W239),
    .Z(W240)
  );

  OR C241 (
    .A(e_input[120]),
    .B(W240),
    .Z(W241)
  );

  OR C242 (
    .A(g_input[121]),
    .B(W241),
    .Z(W242)
  );

  OR C243 (
    .A(e_input[121]),
    .B(W242),
    .Z(W243)
  );

  OR C244 (
    .A(g_input[122]),
    .B(W243),
    .Z(W244)
  );

  OR C245 (
    .A(e_input[122]),
    .B(W244),
    .Z(W245)
  );

  OR C246 (
    .A(g_input[123]),
    .B(W245),
    .Z(W246)
  );

  OR C247 (
    .A(e_input[123]),
    .B(W246),
    .Z(W247)
  );

  OR C248 (
    .A(g_input[124]),
    .B(W247),
    .Z(W248)
  );

  OR C249 (
    .A(e_input[124]),
    .B(W248),
    .Z(W249)
  );

  OR C250 (
    .A(g_input[125]),
    .B(W249),
    .Z(W250)
  );

  OR C251 (
    .A(e_input[125]),
    .B(W250),
    .Z(W251)
  );

  OR C252 (
    .A(g_input[126]),
    .B(W251),
    .Z(W252)
  );

  OR C253 (
    .A(e_input[126]),
    .B(W252),
    .Z(W253)
  );

  OR C254 (
    .A(g_input[127]),
    .B(W253),
    .Z(W254)
  );

  OR C255 (
    .A(e_input[127]),
    .B(W254),
    .Z(W255)
  );

  OR C256 (
    .A(g_input[128]),
    .B(W255),
    .Z(W256)
  );

  OR C257 (
    .A(e_input[128]),
    .B(W256),
    .Z(W257)
  );

  OR C258 (
    .A(g_input[129]),
    .B(W257),
    .Z(W258)
  );

  OR C259 (
    .A(e_input[129]),
    .B(W258),
    .Z(W259)
  );

  OR C260 (
    .A(g_input[130]),
    .B(W259),
    .Z(W260)
  );

  OR C261 (
    .A(e_input[130]),
    .B(W260),
    .Z(W261)
  );

  OR C262 (
    .A(g_input[131]),
    .B(W261),
    .Z(W262)
  );

  OR C263 (
    .A(e_input[131]),
    .B(W262),
    .Z(W263)
  );

  OR C264 (
    .A(g_input[132]),
    .B(W263),
    .Z(W264)
  );

  OR C265 (
    .A(e_input[132]),
    .B(W264),
    .Z(W265)
  );

  OR C266 (
    .A(g_input[133]),
    .B(W265),
    .Z(W266)
  );

  OR C267 (
    .A(e_input[133]),
    .B(W266),
    .Z(W267)
  );

  OR C268 (
    .A(g_input[134]),
    .B(W267),
    .Z(W268)
  );

  OR C269 (
    .A(e_input[134]),
    .B(W268),
    .Z(W269)
  );

  OR C270 (
    .A(g_input[135]),
    .B(W269),
    .Z(W270)
  );

  OR C271 (
    .A(e_input[135]),
    .B(W270),
    .Z(W271)
  );

  OR C272 (
    .A(g_input[136]),
    .B(W271),
    .Z(W272)
  );

  OR C273 (
    .A(e_input[136]),
    .B(W272),
    .Z(W273)
  );

  OR C274 (
    .A(g_input[137]),
    .B(W273),
    .Z(W274)
  );

  OR C275 (
    .A(e_input[137]),
    .B(W274),
    .Z(W275)
  );

  OR C276 (
    .A(g_input[138]),
    .B(W275),
    .Z(W276)
  );

  OR C277 (
    .A(e_input[138]),
    .B(W276),
    .Z(W277)
  );

  OR C278 (
    .A(g_input[139]),
    .B(W277),
    .Z(W278)
  );

  OR C279 (
    .A(e_input[139]),
    .B(W278),
    .Z(W279)
  );

  OR C280 (
    .A(g_input[140]),
    .B(W279),
    .Z(W280)
  );

  OR C281 (
    .A(e_input[140]),
    .B(W280),
    .Z(W281)
  );

  OR C282 (
    .A(g_input[141]),
    .B(W281),
    .Z(W282)
  );

  OR C283 (
    .A(e_input[141]),
    .B(W282),
    .Z(W283)
  );

  OR C284 (
    .A(g_input[142]),
    .B(W283),
    .Z(W284)
  );

  OR C285 (
    .A(e_input[142]),
    .B(W284),
    .Z(W285)
  );

  OR C286 (
    .A(g_input[143]),
    .B(W285),
    .Z(W286)
  );

  OR C287 (
    .A(e_input[143]),
    .B(W286),
    .Z(W287)
  );

  OR C288 (
    .A(g_input[144]),
    .B(W287),
    .Z(W288)
  );

  OR C289 (
    .A(e_input[144]),
    .B(W288),
    .Z(W289)
  );

  OR C290 (
    .A(g_input[145]),
    .B(W289),
    .Z(W290)
  );

  OR C291 (
    .A(e_input[145]),
    .B(W290),
    .Z(W291)
  );

  OR C292 (
    .A(g_input[146]),
    .B(W291),
    .Z(W292)
  );

  OR C293 (
    .A(e_input[146]),
    .B(W292),
    .Z(W293)
  );

  OR C294 (
    .A(g_input[147]),
    .B(W293),
    .Z(W294)
  );

  OR C295 (
    .A(e_input[147]),
    .B(W294),
    .Z(W295)
  );

  OR C296 (
    .A(g_input[148]),
    .B(W295),
    .Z(W296)
  );

  OR C297 (
    .A(e_input[148]),
    .B(W296),
    .Z(W297)
  );

  OR C298 (
    .A(g_input[149]),
    .B(W297),
    .Z(W298)
  );

  OR C299 (
    .A(e_input[149]),
    .B(W298),
    .Z(W299)
  );

  OR C300 (
    .A(g_input[150]),
    .B(W299),
    .Z(W300)
  );

  OR C301 (
    .A(e_input[150]),
    .B(W300),
    .Z(W301)
  );

  OR C302 (
    .A(g_input[151]),
    .B(W301),
    .Z(W302)
  );

  OR C303 (
    .A(e_input[151]),
    .B(W302),
    .Z(W303)
  );

  OR C304 (
    .A(g_input[152]),
    .B(W303),
    .Z(W304)
  );

  OR C305 (
    .A(e_input[152]),
    .B(W304),
    .Z(W305)
  );

  OR C306 (
    .A(g_input[153]),
    .B(W305),
    .Z(W306)
  );

  OR C307 (
    .A(e_input[153]),
    .B(W306),
    .Z(W307)
  );

  OR C308 (
    .A(g_input[154]),
    .B(W307),
    .Z(W308)
  );

  OR C309 (
    .A(e_input[154]),
    .B(W308),
    .Z(W309)
  );

  OR C310 (
    .A(g_input[155]),
    .B(W309),
    .Z(W310)
  );

  OR C311 (
    .A(e_input[155]),
    .B(W310),
    .Z(W311)
  );

  OR C312 (
    .A(g_input[156]),
    .B(W311),
    .Z(W312)
  );

  OR C313 (
    .A(e_input[156]),
    .B(W312),
    .Z(W313)
  );

  OR C314 (
    .A(g_input[157]),
    .B(W313),
    .Z(W314)
  );

  OR C315 (
    .A(e_input[157]),
    .B(W314),
    .Z(W315)
  );

  OR C316 (
    .A(g_input[158]),
    .B(W315),
    .Z(W316)
  );

  OR C317 (
    .A(e_input[158]),
    .B(W316),
    .Z(W317)
  );

  OR C318 (
    .A(g_input[159]),
    .B(W317),
    .Z(W318)
  );

  OR C319 (
    .A(e_input[159]),
    .B(W318),
    .Z(W319)
  );

  OR C320 (
    .A(g_input[160]),
    .B(W319),
    .Z(W320)
  );

  OR C321 (
    .A(e_input[160]),
    .B(W320),
    .Z(W321)
  );

  OR C322 (
    .A(g_input[161]),
    .B(W321),
    .Z(W322)
  );

  OR C323 (
    .A(e_input[161]),
    .B(W322),
    .Z(W323)
  );

  OR C324 (
    .A(g_input[162]),
    .B(W323),
    .Z(W324)
  );

  OR C325 (
    .A(e_input[162]),
    .B(W324),
    .Z(W325)
  );

  OR C326 (
    .A(g_input[163]),
    .B(W325),
    .Z(W326)
  );

  OR C327 (
    .A(e_input[163]),
    .B(W326),
    .Z(W327)
  );

  OR C328 (
    .A(g_input[164]),
    .B(W327),
    .Z(W328)
  );

  OR C329 (
    .A(e_input[164]),
    .B(W328),
    .Z(W329)
  );

  OR C330 (
    .A(g_input[165]),
    .B(W329),
    .Z(W330)
  );

  OR C331 (
    .A(e_input[165]),
    .B(W330),
    .Z(W331)
  );

  OR C332 (
    .A(g_input[166]),
    .B(W331),
    .Z(W332)
  );

  OR C333 (
    .A(e_input[166]),
    .B(W332),
    .Z(W333)
  );

  OR C334 (
    .A(g_input[167]),
    .B(W333),
    .Z(W334)
  );

  OR C335 (
    .A(e_input[167]),
    .B(W334),
    .Z(W335)
  );

  OR C336 (
    .A(g_input[168]),
    .B(W335),
    .Z(W336)
  );

  OR C337 (
    .A(e_input[168]),
    .B(W336),
    .Z(W337)
  );

  OR C338 (
    .A(g_input[169]),
    .B(W337),
    .Z(W338)
  );

  OR C339 (
    .A(e_input[169]),
    .B(W338),
    .Z(W339)
  );

  OR C340 (
    .A(g_input[170]),
    .B(W339),
    .Z(W340)
  );

  OR C341 (
    .A(e_input[170]),
    .B(W340),
    .Z(W341)
  );

  OR C342 (
    .A(g_input[171]),
    .B(W341),
    .Z(W342)
  );

  OR C343 (
    .A(e_input[171]),
    .B(W342),
    .Z(W343)
  );

  OR C344 (
    .A(g_input[172]),
    .B(W343),
    .Z(W344)
  );

  OR C345 (
    .A(e_input[172]),
    .B(W344),
    .Z(W345)
  );

  OR C346 (
    .A(g_input[173]),
    .B(W345),
    .Z(W346)
  );

  OR C347 (
    .A(e_input[173]),
    .B(W346),
    .Z(W347)
  );

  OR C348 (
    .A(g_input[174]),
    .B(W347),
    .Z(W348)
  );

  OR C349 (
    .A(e_input[174]),
    .B(W348),
    .Z(W349)
  );

  OR C350 (
    .A(g_input[175]),
    .B(W349),
    .Z(W350)
  );

  OR C351 (
    .A(e_input[175]),
    .B(W350),
    .Z(W351)
  );

  OR C352 (
    .A(g_input[176]),
    .B(W351),
    .Z(W352)
  );

  OR C353 (
    .A(e_input[176]),
    .B(W352),
    .Z(W353)
  );

  OR C354 (
    .A(g_input[177]),
    .B(W353),
    .Z(W354)
  );

  OR C355 (
    .A(e_input[177]),
    .B(W354),
    .Z(W355)
  );

  OR C356 (
    .A(g_input[178]),
    .B(W355),
    .Z(W356)
  );

  OR C357 (
    .A(e_input[178]),
    .B(W356),
    .Z(W357)
  );

  OR C358 (
    .A(g_input[179]),
    .B(W357),
    .Z(W358)
  );

  OR C359 (
    .A(e_input[179]),
    .B(W358),
    .Z(W359)
  );

  OR C360 (
    .A(g_input[180]),
    .B(W359),
    .Z(W360)
  );

  OR C361 (
    .A(e_input[180]),
    .B(W360),
    .Z(W361)
  );

  OR C362 (
    .A(g_input[181]),
    .B(W361),
    .Z(W362)
  );

  OR C363 (
    .A(e_input[181]),
    .B(W362),
    .Z(W363)
  );

  OR C364 (
    .A(g_input[182]),
    .B(W363),
    .Z(W364)
  );

  OR C365 (
    .A(e_input[182]),
    .B(W364),
    .Z(W365)
  );

  OR C366 (
    .A(g_input[183]),
    .B(W365),
    .Z(W366)
  );

  OR C367 (
    .A(e_input[183]),
    .B(W366),
    .Z(W367)
  );

  OR C368 (
    .A(g_input[184]),
    .B(W367),
    .Z(W368)
  );

  OR C369 (
    .A(e_input[184]),
    .B(W368),
    .Z(W369)
  );

  OR C370 (
    .A(g_input[185]),
    .B(W369),
    .Z(W370)
  );

  OR C371 (
    .A(e_input[185]),
    .B(W370),
    .Z(W371)
  );

  OR C372 (
    .A(g_input[186]),
    .B(W371),
    .Z(W372)
  );

  OR C373 (
    .A(e_input[186]),
    .B(W372),
    .Z(W373)
  );

  OR C374 (
    .A(g_input[187]),
    .B(W373),
    .Z(W374)
  );

  OR C375 (
    .A(e_input[187]),
    .B(W374),
    .Z(W375)
  );

  OR C376 (
    .A(g_input[188]),
    .B(W375),
    .Z(W376)
  );

  OR C377 (
    .A(e_input[188]),
    .B(W376),
    .Z(W377)
  );

  OR C378 (
    .A(g_input[189]),
    .B(W377),
    .Z(W378)
  );

  OR C379 (
    .A(e_input[189]),
    .B(W378),
    .Z(W379)
  );

  OR C380 (
    .A(g_input[190]),
    .B(W379),
    .Z(W380)
  );

  OR C381 (
    .A(e_input[190]),
    .B(W380),
    .Z(W381)
  );

  OR C382 (
    .A(g_input[191]),
    .B(W381),
    .Z(W382)
  );

  OR C383 (
    .A(e_input[191]),
    .B(W382),
    .Z(W383)
  );

  OR C384 (
    .A(g_input[192]),
    .B(W383),
    .Z(W384)
  );

  OR C385 (
    .A(e_input[192]),
    .B(W384),
    .Z(W385)
  );

  OR C386 (
    .A(g_input[193]),
    .B(W385),
    .Z(W386)
  );

  OR C387 (
    .A(e_input[193]),
    .B(W386),
    .Z(W387)
  );

  OR C388 (
    .A(g_input[194]),
    .B(W387),
    .Z(W388)
  );

  OR C389 (
    .A(e_input[194]),
    .B(W388),
    .Z(W389)
  );

  OR C390 (
    .A(g_input[195]),
    .B(W389),
    .Z(W390)
  );

  OR C391 (
    .A(e_input[195]),
    .B(W390),
    .Z(W391)
  );

  OR C392 (
    .A(g_input[196]),
    .B(W391),
    .Z(W392)
  );

  OR C393 (
    .A(e_input[196]),
    .B(W392),
    .Z(W393)
  );

  OR C394 (
    .A(g_input[197]),
    .B(W393),
    .Z(W394)
  );

  OR C395 (
    .A(e_input[197]),
    .B(W394),
    .Z(W395)
  );

  OR C396 (
    .A(g_input[198]),
    .B(W395),
    .Z(W396)
  );

  OR C397 (
    .A(e_input[198]),
    .B(W396),
    .Z(W397)
  );

  OR C398 (
    .A(g_input[199]),
    .B(W397),
    .Z(W398)
  );

  OR C399 (
    .A(e_input[199]),
    .B(W398),
    .Z(W399)
  );

  OR C400 (
    .A(g_input[200]),
    .B(W399),
    .Z(W400)
  );

  OR C401 (
    .A(e_input[200]),
    .B(W400),
    .Z(W401)
  );

  OR C402 (
    .A(g_input[201]),
    .B(W401),
    .Z(W402)
  );

  OR C403 (
    .A(e_input[201]),
    .B(W402),
    .Z(W403)
  );

  OR C404 (
    .A(g_input[202]),
    .B(W403),
    .Z(W404)
  );

  OR C405 (
    .A(e_input[202]),
    .B(W404),
    .Z(W405)
  );

  OR C406 (
    .A(g_input[203]),
    .B(W405),
    .Z(W406)
  );

  OR C407 (
    .A(e_input[203]),
    .B(W406),
    .Z(W407)
  );

  OR C408 (
    .A(g_input[204]),
    .B(W407),
    .Z(W408)
  );

  OR C409 (
    .A(e_input[204]),
    .B(W408),
    .Z(W409)
  );

  OR C410 (
    .A(g_input[205]),
    .B(W409),
    .Z(W410)
  );

  OR C411 (
    .A(e_input[205]),
    .B(W410),
    .Z(W411)
  );

  OR C412 (
    .A(g_input[206]),
    .B(W411),
    .Z(W412)
  );

  OR C413 (
    .A(e_input[206]),
    .B(W412),
    .Z(W413)
  );

  OR C414 (
    .A(g_input[207]),
    .B(W413),
    .Z(W414)
  );

  OR C415 (
    .A(e_input[207]),
    .B(W414),
    .Z(W415)
  );

  OR C416 (
    .A(g_input[208]),
    .B(W415),
    .Z(W416)
  );

  OR C417 (
    .A(e_input[208]),
    .B(W416),
    .Z(W417)
  );

  OR C418 (
    .A(g_input[209]),
    .B(W417),
    .Z(W418)
  );

  OR C419 (
    .A(e_input[209]),
    .B(W418),
    .Z(W419)
  );

  OR C420 (
    .A(g_input[210]),
    .B(W419),
    .Z(W420)
  );

  OR C421 (
    .A(e_input[210]),
    .B(W420),
    .Z(W421)
  );

  OR C422 (
    .A(g_input[211]),
    .B(W421),
    .Z(W422)
  );

  OR C423 (
    .A(e_input[211]),
    .B(W422),
    .Z(W423)
  );

  OR C424 (
    .A(g_input[212]),
    .B(W423),
    .Z(W424)
  );

  OR C425 (
    .A(e_input[212]),
    .B(W424),
    .Z(W425)
  );

  OR C426 (
    .A(g_input[213]),
    .B(W425),
    .Z(W426)
  );

  OR C427 (
    .A(e_input[213]),
    .B(W426),
    .Z(W427)
  );

  OR C428 (
    .A(g_input[214]),
    .B(W427),
    .Z(W428)
  );

  OR C429 (
    .A(e_input[214]),
    .B(W428),
    .Z(W429)
  );

  OR C430 (
    .A(g_input[215]),
    .B(W429),
    .Z(W430)
  );

  OR C431 (
    .A(e_input[215]),
    .B(W430),
    .Z(W431)
  );

  OR C432 (
    .A(g_input[216]),
    .B(W431),
    .Z(W432)
  );

  OR C433 (
    .A(e_input[216]),
    .B(W432),
    .Z(W433)
  );

  OR C434 (
    .A(g_input[217]),
    .B(W433),
    .Z(W434)
  );

  OR C435 (
    .A(e_input[217]),
    .B(W434),
    .Z(W435)
  );

  OR C436 (
    .A(g_input[218]),
    .B(W435),
    .Z(W436)
  );

  OR C437 (
    .A(e_input[218]),
    .B(W436),
    .Z(W437)
  );

  OR C438 (
    .A(g_input[219]),
    .B(W437),
    .Z(W438)
  );

  OR C439 (
    .A(e_input[219]),
    .B(W438),
    .Z(W439)
  );

  OR C440 (
    .A(g_input[220]),
    .B(W439),
    .Z(W440)
  );

  OR C441 (
    .A(e_input[220]),
    .B(W440),
    .Z(W441)
  );

  OR C442 (
    .A(g_input[221]),
    .B(W441),
    .Z(W442)
  );

  OR C443 (
    .A(e_input[221]),
    .B(W442),
    .Z(W443)
  );

  OR C444 (
    .A(g_input[222]),
    .B(W443),
    .Z(W444)
  );

  OR C445 (
    .A(e_input[222]),
    .B(W444),
    .Z(W445)
  );

  OR C446 (
    .A(g_input[223]),
    .B(W445),
    .Z(W446)
  );

  OR C447 (
    .A(e_input[223]),
    .B(W446),
    .Z(W447)
  );

  OR C448 (
    .A(g_input[224]),
    .B(W447),
    .Z(W448)
  );

  OR C449 (
    .A(e_input[224]),
    .B(W448),
    .Z(W449)
  );

  OR C450 (
    .A(g_input[225]),
    .B(W449),
    .Z(W450)
  );

  OR C451 (
    .A(e_input[225]),
    .B(W450),
    .Z(W451)
  );

  OR C452 (
    .A(g_input[226]),
    .B(W451),
    .Z(W452)
  );

  OR C453 (
    .A(e_input[226]),
    .B(W452),
    .Z(W453)
  );

  OR C454 (
    .A(g_input[227]),
    .B(W453),
    .Z(W454)
  );

  OR C455 (
    .A(e_input[227]),
    .B(W454),
    .Z(W455)
  );

  OR C456 (
    .A(g_input[228]),
    .B(W455),
    .Z(W456)
  );

  OR C457 (
    .A(e_input[228]),
    .B(W456),
    .Z(W457)
  );

  OR C458 (
    .A(g_input[229]),
    .B(W457),
    .Z(W458)
  );

  OR C459 (
    .A(e_input[229]),
    .B(W458),
    .Z(W459)
  );

  OR C460 (
    .A(g_input[230]),
    .B(W459),
    .Z(W460)
  );

  OR C461 (
    .A(e_input[230]),
    .B(W460),
    .Z(W461)
  );

  OR C462 (
    .A(g_input[231]),
    .B(W461),
    .Z(W462)
  );

  OR C463 (
    .A(e_input[231]),
    .B(W462),
    .Z(W463)
  );

  OR C464 (
    .A(g_input[232]),
    .B(W463),
    .Z(W464)
  );

  OR C465 (
    .A(e_input[232]),
    .B(W464),
    .Z(W465)
  );

  OR C466 (
    .A(g_input[233]),
    .B(W465),
    .Z(W466)
  );

  OR C467 (
    .A(e_input[233]),
    .B(W466),
    .Z(W467)
  );

  OR C468 (
    .A(g_input[234]),
    .B(W467),
    .Z(W468)
  );

  OR C469 (
    .A(e_input[234]),
    .B(W468),
    .Z(W469)
  );

  OR C470 (
    .A(g_input[235]),
    .B(W469),
    .Z(W470)
  );

  OR C471 (
    .A(e_input[235]),
    .B(W470),
    .Z(W471)
  );

  OR C472 (
    .A(g_input[236]),
    .B(W471),
    .Z(W472)
  );

  OR C473 (
    .A(e_input[236]),
    .B(W472),
    .Z(W473)
  );

  OR C474 (
    .A(g_input[237]),
    .B(W473),
    .Z(W474)
  );

  OR C475 (
    .A(e_input[237]),
    .B(W474),
    .Z(W475)
  );

  OR C476 (
    .A(g_input[238]),
    .B(W475),
    .Z(W476)
  );

  OR C477 (
    .A(e_input[238]),
    .B(W476),
    .Z(W477)
  );

  OR C478 (
    .A(g_input[239]),
    .B(W477),
    .Z(W478)
  );

  OR C479 (
    .A(e_input[239]),
    .B(W478),
    .Z(W479)
  );

  OR C480 (
    .A(g_input[240]),
    .B(W479),
    .Z(W480)
  );

  OR C481 (
    .A(e_input[240]),
    .B(W480),
    .Z(W481)
  );

  OR C482 (
    .A(g_input[241]),
    .B(W481),
    .Z(W482)
  );

  OR C483 (
    .A(e_input[241]),
    .B(W482),
    .Z(W483)
  );

  OR C484 (
    .A(g_input[242]),
    .B(W483),
    .Z(W484)
  );

  OR C485 (
    .A(e_input[242]),
    .B(W484),
    .Z(W485)
  );

  OR C486 (
    .A(g_input[243]),
    .B(W485),
    .Z(W486)
  );

  OR C487 (
    .A(e_input[243]),
    .B(W486),
    .Z(W487)
  );

  OR C488 (
    .A(g_input[244]),
    .B(W487),
    .Z(W488)
  );

  OR C489 (
    .A(e_input[244]),
    .B(W488),
    .Z(W489)
  );

  OR C490 (
    .A(g_input[245]),
    .B(W489),
    .Z(W490)
  );

  OR C491 (
    .A(e_input[245]),
    .B(W490),
    .Z(W491)
  );

  OR C492 (
    .A(g_input[246]),
    .B(W491),
    .Z(W492)
  );

  OR C493 (
    .A(e_input[246]),
    .B(W492),
    .Z(W493)
  );

  OR C494 (
    .A(g_input[247]),
    .B(W493),
    .Z(W494)
  );

  OR C495 (
    .A(e_input[247]),
    .B(W494),
    .Z(W495)
  );

  OR C496 (
    .A(g_input[248]),
    .B(W495),
    .Z(W496)
  );

  OR C497 (
    .A(e_input[248]),
    .B(W496),
    .Z(W497)
  );

  OR C498 (
    .A(g_input[249]),
    .B(W497),
    .Z(W498)
  );

  OR C499 (
    .A(e_input[249]),
    .B(W498),
    .Z(W499)
  );

  OR C500 (
    .A(g_input[250]),
    .B(W499),
    .Z(W500)
  );

  OR C501 (
    .A(e_input[250]),
    .B(W500),
    .Z(W501)
  );

  OR C502 (
    .A(g_input[251]),
    .B(W501),
    .Z(W502)
  );

  OR C503 (
    .A(e_input[251]),
    .B(W502),
    .Z(W503)
  );

  OR C504 (
    .A(g_input[252]),
    .B(W503),
    .Z(W504)
  );

  OR C505 (
    .A(e_input[252]),
    .B(W504),
    .Z(W505)
  );

  OR C506 (
    .A(g_input[253]),
    .B(W505),
    .Z(W506)
  );

  OR C507 (
    .A(e_input[253]),
    .B(W506),
    .Z(W507)
  );

  OR C508 (
    .A(g_input[254]),
    .B(W507),
    .Z(W508)
  );

  OR C509 (
    .A(e_input[254]),
    .B(W508),
    .Z(W509)
  );

  OR C510 (
    .A(g_input[255]),
    .B(W509),
    .Z(W510)
  );

  OR C511 (
    .A(e_input[255]),
    .B(W510),
    .Z(o)
  );
endmodule
